package ram_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "ram_txn.sv"
  `include "ram_sequencer.sv"
  `include "ram_driver.sv"
  `include "ram_monitor.sv"
  `include "ram_agent.sv"
  `include "ram_env.sv"
  `include "ram_test.sv"
endpackage
